
module soc_system (
	button_pio_external_connection_export,
	clk_clk,
	ctrl_out_export,
	dipsw_pio_external_connection_export,
	hps_0_f2h_cold_reset_req_reset_n,
	hps_0_f2h_debug_reset_req_reset_n,
	hps_0_f2h_stm_hw_events_stm_hwevents,
	hps_0_f2h_warm_reset_req_reset_n,
	hps_0_h2f_reset_reset_n,
	hps_0_hps_io_hps_io_emac1_inst_TX_CLK,
	hps_0_hps_io_hps_io_emac1_inst_TXD0,
	hps_0_hps_io_hps_io_emac1_inst_TXD1,
	hps_0_hps_io_hps_io_emac1_inst_TXD2,
	hps_0_hps_io_hps_io_emac1_inst_TXD3,
	hps_0_hps_io_hps_io_emac1_inst_RXD0,
	hps_0_hps_io_hps_io_emac1_inst_MDIO,
	hps_0_hps_io_hps_io_emac1_inst_MDC,
	hps_0_hps_io_hps_io_emac1_inst_RX_CTL,
	hps_0_hps_io_hps_io_emac1_inst_TX_CTL,
	hps_0_hps_io_hps_io_emac1_inst_RX_CLK,
	hps_0_hps_io_hps_io_emac1_inst_RXD1,
	hps_0_hps_io_hps_io_emac1_inst_RXD2,
	hps_0_hps_io_hps_io_emac1_inst_RXD3,
	hps_0_hps_io_hps_io_sdio_inst_CMD,
	hps_0_hps_io_hps_io_sdio_inst_D0,
	hps_0_hps_io_hps_io_sdio_inst_D1,
	hps_0_hps_io_hps_io_sdio_inst_CLK,
	hps_0_hps_io_hps_io_sdio_inst_D2,
	hps_0_hps_io_hps_io_sdio_inst_D3,
	hps_0_hps_io_hps_io_usb1_inst_D0,
	hps_0_hps_io_hps_io_usb1_inst_D1,
	hps_0_hps_io_hps_io_usb1_inst_D2,
	hps_0_hps_io_hps_io_usb1_inst_D3,
	hps_0_hps_io_hps_io_usb1_inst_D4,
	hps_0_hps_io_hps_io_usb1_inst_D5,
	hps_0_hps_io_hps_io_usb1_inst_D6,
	hps_0_hps_io_hps_io_usb1_inst_D7,
	hps_0_hps_io_hps_io_usb1_inst_CLK,
	hps_0_hps_io_hps_io_usb1_inst_STP,
	hps_0_hps_io_hps_io_usb1_inst_DIR,
	hps_0_hps_io_hps_io_usb1_inst_NXT,
	hps_0_hps_io_hps_io_spim1_inst_CLK,
	hps_0_hps_io_hps_io_spim1_inst_MOSI,
	hps_0_hps_io_hps_io_spim1_inst_MISO,
	hps_0_hps_io_hps_io_spim1_inst_SS0,
	hps_0_hps_io_hps_io_uart0_inst_RX,
	hps_0_hps_io_hps_io_uart0_inst_TX,
	hps_0_hps_io_hps_io_i2c0_inst_SDA,
	hps_0_hps_io_hps_io_i2c0_inst_SCL,
	hps_0_hps_io_hps_io_i2c1_inst_SDA,
	hps_0_hps_io_hps_io_i2c1_inst_SCL,
	hps_0_hps_io_hps_io_gpio_inst_GPIO09,
	hps_0_hps_io_hps_io_gpio_inst_GPIO35,
	hps_0_hps_io_hps_io_gpio_inst_GPIO40,
	hps_0_hps_io_hps_io_gpio_inst_GPIO53,
	hps_0_hps_io_hps_io_gpio_inst_GPIO54,
	hps_0_hps_io_hps_io_gpio_inst_GPIO61,
	i2c_ext_sda_in,
	i2c_ext_scl_in,
	i2c_ext_sda_oe,
	i2c_ext_scl_oe,
	i2c_ext_1_sda_in,
	i2c_ext_1_scl_in,
	i2c_ext_1_sda_oe,
	i2c_ext_1_scl_oe,
	i2c_int_sda_in,
	i2c_int_scl_in,
	i2c_int_sda_oe,
	i2c_int_scl_oe,
	led_pio_external_connection_export,
	memory_mem_a,
	memory_mem_ba,
	memory_mem_ck,
	memory_mem_ck_n,
	memory_mem_cke,
	memory_mem_cs_n,
	memory_mem_ras_n,
	memory_mem_cas_n,
	memory_mem_we_n,
	memory_mem_reset_n,
	memory_mem_dq,
	memory_mem_dqs,
	memory_mem_dqs_n,
	memory_mem_odt,
	memory_mem_dm,
	memory_oct_rzqin,
	pulse_gpio_pio_external_connection_export,
	pulse_length_ch2_para_export,
	pulse_length_ch3_para_export,
	pulse_length_ch4_para_export,
	pulse_length_para_export,
	pulse_length_pio_0_external_connection_export,
	pulse_length_pio_10_external_connection_export,
	pulse_length_pio_11_external_connection_export,
	pulse_length_pio_12_external_connection_export,
	pulse_length_pio_13_external_connection_export,
	pulse_length_pio_14_external_connection_export,
	pulse_length_pio_15_external_connection_export,
	pulse_length_pio_16_external_connection_export,
	pulse_length_pio_17_external_connection_export,
	pulse_length_pio_18_external_connection_export,
	pulse_length_pio_19_external_connection_export,
	pulse_length_pio_1_external_connection_export,
	pulse_length_pio_20_external_connection_export,
	pulse_length_pio_21_external_connection_export,
	pulse_length_pio_22_external_connection_export,
	pulse_length_pio_23_external_connection_export,
	pulse_length_pio_24_external_connection_export,
	pulse_length_pio_25_external_connection_export,
	pulse_length_pio_26_external_connection_export,
	pulse_length_pio_27_external_connection_export,
	pulse_length_pio_28_external_connection_export,
	pulse_length_pio_29_external_connection_export,
	pulse_length_pio_2_external_connection_export,
	pulse_length_pio_30_external_connection_export,
	pulse_length_pio_31_external_connection_export,
	pulse_length_pio_32_external_connection_export,
	pulse_length_pio_33_external_connection_export,
	pulse_length_pio_34_external_connection_export,
	pulse_length_pio_35_external_connection_export,
	pulse_length_pio_3_external_connection_export,
	pulse_length_pio_4_external_connection_export,
	pulse_length_pio_5_external_connection_export,
	pulse_length_pio_6_external_connection_export,
	pulse_length_pio_7_external_connection_export,
	pulse_length_pio_8_external_connection_export,
	pulse_length_pio_9_external_connection_export,
	reset_reset_n);	

	input	[1:0]	button_pio_external_connection_export;
	input		clk_clk;
	output	[31:0]	ctrl_out_export;
	input	[3:0]	dipsw_pio_external_connection_export;
	input		hps_0_f2h_cold_reset_req_reset_n;
	input		hps_0_f2h_debug_reset_req_reset_n;
	input	[27:0]	hps_0_f2h_stm_hw_events_stm_hwevents;
	input		hps_0_f2h_warm_reset_req_reset_n;
	output		hps_0_h2f_reset_reset_n;
	output		hps_0_hps_io_hps_io_emac1_inst_TX_CLK;
	output		hps_0_hps_io_hps_io_emac1_inst_TXD0;
	output		hps_0_hps_io_hps_io_emac1_inst_TXD1;
	output		hps_0_hps_io_hps_io_emac1_inst_TXD2;
	output		hps_0_hps_io_hps_io_emac1_inst_TXD3;
	input		hps_0_hps_io_hps_io_emac1_inst_RXD0;
	inout		hps_0_hps_io_hps_io_emac1_inst_MDIO;
	output		hps_0_hps_io_hps_io_emac1_inst_MDC;
	input		hps_0_hps_io_hps_io_emac1_inst_RX_CTL;
	output		hps_0_hps_io_hps_io_emac1_inst_TX_CTL;
	input		hps_0_hps_io_hps_io_emac1_inst_RX_CLK;
	input		hps_0_hps_io_hps_io_emac1_inst_RXD1;
	input		hps_0_hps_io_hps_io_emac1_inst_RXD2;
	input		hps_0_hps_io_hps_io_emac1_inst_RXD3;
	inout		hps_0_hps_io_hps_io_sdio_inst_CMD;
	inout		hps_0_hps_io_hps_io_sdio_inst_D0;
	inout		hps_0_hps_io_hps_io_sdio_inst_D1;
	output		hps_0_hps_io_hps_io_sdio_inst_CLK;
	inout		hps_0_hps_io_hps_io_sdio_inst_D2;
	inout		hps_0_hps_io_hps_io_sdio_inst_D3;
	inout		hps_0_hps_io_hps_io_usb1_inst_D0;
	inout		hps_0_hps_io_hps_io_usb1_inst_D1;
	inout		hps_0_hps_io_hps_io_usb1_inst_D2;
	inout		hps_0_hps_io_hps_io_usb1_inst_D3;
	inout		hps_0_hps_io_hps_io_usb1_inst_D4;
	inout		hps_0_hps_io_hps_io_usb1_inst_D5;
	inout		hps_0_hps_io_hps_io_usb1_inst_D6;
	inout		hps_0_hps_io_hps_io_usb1_inst_D7;
	input		hps_0_hps_io_hps_io_usb1_inst_CLK;
	output		hps_0_hps_io_hps_io_usb1_inst_STP;
	input		hps_0_hps_io_hps_io_usb1_inst_DIR;
	input		hps_0_hps_io_hps_io_usb1_inst_NXT;
	output		hps_0_hps_io_hps_io_spim1_inst_CLK;
	output		hps_0_hps_io_hps_io_spim1_inst_MOSI;
	input		hps_0_hps_io_hps_io_spim1_inst_MISO;
	output		hps_0_hps_io_hps_io_spim1_inst_SS0;
	input		hps_0_hps_io_hps_io_uart0_inst_RX;
	output		hps_0_hps_io_hps_io_uart0_inst_TX;
	inout		hps_0_hps_io_hps_io_i2c0_inst_SDA;
	inout		hps_0_hps_io_hps_io_i2c0_inst_SCL;
	inout		hps_0_hps_io_hps_io_i2c1_inst_SDA;
	inout		hps_0_hps_io_hps_io_i2c1_inst_SCL;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO09;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO35;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO40;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO53;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO54;
	inout		hps_0_hps_io_hps_io_gpio_inst_GPIO61;
	input		i2c_ext_sda_in;
	input		i2c_ext_scl_in;
	output		i2c_ext_sda_oe;
	output		i2c_ext_scl_oe;
	input		i2c_ext_1_sda_in;
	input		i2c_ext_1_scl_in;
	output		i2c_ext_1_sda_oe;
	output		i2c_ext_1_scl_oe;
	input		i2c_int_sda_in;
	input		i2c_int_scl_in;
	output		i2c_int_sda_oe;
	output		i2c_int_scl_oe;
	output	[6:0]	led_pio_external_connection_export;
	output	[14:0]	memory_mem_a;
	output	[2:0]	memory_mem_ba;
	output		memory_mem_ck;
	output		memory_mem_ck_n;
	output		memory_mem_cke;
	output		memory_mem_cs_n;
	output		memory_mem_ras_n;
	output		memory_mem_cas_n;
	output		memory_mem_we_n;
	output		memory_mem_reset_n;
	inout	[31:0]	memory_mem_dq;
	inout	[3:0]	memory_mem_dqs;
	inout	[3:0]	memory_mem_dqs_n;
	output		memory_mem_odt;
	output	[3:0]	memory_mem_dm;
	input		memory_oct_rzqin;
	output	[6:0]	pulse_gpio_pio_external_connection_export;
	output	[31:0]	pulse_length_ch2_para_export;
	output	[31:0]	pulse_length_ch3_para_export;
	output	[31:0]	pulse_length_ch4_para_export;
	output	[31:0]	pulse_length_para_export;
	output	[31:0]	pulse_length_pio_0_external_connection_export;
	output	[31:0]	pulse_length_pio_10_external_connection_export;
	output	[31:0]	pulse_length_pio_11_external_connection_export;
	output	[31:0]	pulse_length_pio_12_external_connection_export;
	output	[31:0]	pulse_length_pio_13_external_connection_export;
	output	[31:0]	pulse_length_pio_14_external_connection_export;
	output	[31:0]	pulse_length_pio_15_external_connection_export;
	output	[31:0]	pulse_length_pio_16_external_connection_export;
	output	[31:0]	pulse_length_pio_17_external_connection_export;
	output	[31:0]	pulse_length_pio_18_external_connection_export;
	output	[31:0]	pulse_length_pio_19_external_connection_export;
	output	[31:0]	pulse_length_pio_1_external_connection_export;
	output	[31:0]	pulse_length_pio_20_external_connection_export;
	output	[31:0]	pulse_length_pio_21_external_connection_export;
	output	[31:0]	pulse_length_pio_22_external_connection_export;
	output	[31:0]	pulse_length_pio_23_external_connection_export;
	output	[31:0]	pulse_length_pio_24_external_connection_export;
	output	[31:0]	pulse_length_pio_25_external_connection_export;
	output	[31:0]	pulse_length_pio_26_external_connection_export;
	output	[31:0]	pulse_length_pio_27_external_connection_export;
	output	[31:0]	pulse_length_pio_28_external_connection_export;
	output	[31:0]	pulse_length_pio_29_external_connection_export;
	output	[31:0]	pulse_length_pio_2_external_connection_export;
	output	[31:0]	pulse_length_pio_30_external_connection_export;
	output	[31:0]	pulse_length_pio_31_external_connection_export;
	output	[31:0]	pulse_length_pio_32_external_connection_export;
	output	[31:0]	pulse_length_pio_33_external_connection_export;
	output	[31:0]	pulse_length_pio_34_external_connection_export;
	output	[31:0]	pulse_length_pio_35_external_connection_export;
	output	[31:0]	pulse_length_pio_3_external_connection_export;
	output	[31:0]	pulse_length_pio_4_external_connection_export;
	output	[31:0]	pulse_length_pio_5_external_connection_export;
	output	[31:0]	pulse_length_pio_6_external_connection_export;
	output	[31:0]	pulse_length_pio_7_external_connection_export;
	output	[31:0]	pulse_length_pio_8_external_connection_export;
	output	[31:0]	pulse_length_pio_9_external_connection_export;
	input		reset_reset_n;
endmodule
